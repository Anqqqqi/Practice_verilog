module sync_fifo #(
parameter DATA_WIDTH = 8, 
arameter DATA_DEPTH = 128)
(
    
);
endmodule